library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;


entity bin2bcd_12bit is  -- Converts binary numbers to a bcd display 
    Port ( binIN : in  STD_LOGIC_VECTOR (10 downto 0); -- the binary number in to be converted
           ones : out  STD_LOGIC_VECTOR (4 downto 0); -- return of the ones in 7 segs
           tens : out  STD_LOGIC_VECTOR (4 downto 0); -- return of the tens in 7 segs
           hundreds : out  STD_LOGIC_VECTOR (4 downto 0); -- return of the hundreds in 7 segs
           thousands : out  STD_LOGIC_VECTOR (4 downto 0) -- return of the thousands in 7 segs
          );
end bin2bcd_12bit;

architecture Behavioral of bin2bcd_12bit is

begin

bcd1: process(binIN)

  -- temporary variable
  variable temp : STD_LOGIC_VECTOR (10 downto 0);
  
  -- variable to store the output BCD number
  -- organized as follows
  -- thousands = bcd(15 downto 12)
  -- hundreds = bcd(11 downto 8)
  -- tens = bcd(7 downto 4)
  -- units = bcd(3 downto 0)
  variable bcd : UNSIGNED (15 downto 0) := (others => '0');

  -- by
  -- https://en.wikipedia.org/wiki/Double_dabble
  
  begin
    -- zero the bcd variable
    bcd := (others => '0');
    
    -- read input into temp variable
    temp(10 downto 0) := binIN;
    
    -- cycle 12 times as we have 12 input bits
    -- this could be optimized, we do not need to check and add 3 for the 
    -- first 3 iterations as the number can never be >4
    for i in 0 to 10 loop
    
      if bcd(3 downto 0) > 4 then 
        bcd(3 downto 0) := bcd(3 downto 0) + 3;
      end if;
      
      if bcd(7 downto 4) > 4 then 
        bcd(7 downto 4) := bcd(7 downto 4) + 3;
      end if;
    
      if bcd(11 downto 8) > 4 then  
        bcd(11 downto 8) := bcd(11 downto 8) + 3;
      end if;
    
      -- thousands can't be >4 for a 12-bit input number
      -- so don't need to do anything to upper 4 bits of bcd
    
      -- shift bcd left by 1 bit, copy MSB of temp into LSB of bcd
      bcd := bcd(14 downto 0) & temp(10);
    
      -- shift temp left by 1 bit
      temp := temp(9 downto 0) & '0';
    
    end loop;
 
    -- set outputs
    ones <= '0' & STD_LOGIC_VECTOR(bcd(3 downto 0));
    tens <= '0' & STD_LOGIC_VECTOR(bcd(7 downto 4));
    hundreds <= '0' & STD_LOGIC_VECTOR(bcd(11 downto 8));
    thousands <= '0' & STD_LOGIC_VECTOR(bcd(15 downto 12));
  
  end process bcd1;            
  
end Behavioral;